package sgls;
 `include "clk_gen.sv"
 `include "rst_gen.sv"
 `include "simulation.sv"
 `include "comparison.sv"
 `include "run.sv"
endpackage
