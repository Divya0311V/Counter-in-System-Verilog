//signals from design
interface counter_sgl;
  logic clk;
  logic rst;
  logic exact;
  logic [7:0]out;
endinterface
